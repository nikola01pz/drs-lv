library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity sevenSegmentBTNU is
	port( 
	);
end sevenSegmentBTNU;

architecture Behavioral of sevenSegmentBTNU is

begin


end Behavioral;

